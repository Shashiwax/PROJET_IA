* RC low-pass filter - first order

.param Rval = {RVAL}
.param Cval = {CVAL}

Vin in 0 AC 1
R1 in out {Rval}
C1 out 0 {Cval}

.ac dec 100 1 1Meg
.meas ac fcut WHEN vdb(out) = -3 CROSS=1

.end
