* RC low-pass filter - first order

* ---------- Paramètres ----------
.param Rval = 1k
.param Cval = 1u

* ---------- Source d'entrée ----------
* Source AC de 1 V efficace
Vin in 0 AC 1

* ---------- Réseau RC ----------
* R entre l'entrée et la sortie
R1 in out {Rval}
* C entre la sortie et la masse
C1 out 0 {Cval}

* ---------- Analyse AC ----------
* Balayage en fréquence : 100 points par décade
* de 1 Hz à 1 MHz
.ac dec 100 1 1Meg

* ---------- Mesure de la fréquence de coupure ----------
* Fréquence pour laquelle le gain en dB sur la sortie vaut -3 dB
.meas ac fcut WHEN vdb(out) = -3 CROSS=1

* (Optionnel) Impression du gain en dB
* .print ac vdb(v(out))

.end
